// ?????????? ?????? RS-???????? ? ??? ??????????: 
module RStrigger (out,x,xdop); 
 
// ??????????? ??????????    
  // ??????? ? ????????: x � S; xdop � R; out - !Q 
   input x,xdop; 
   output out; 
 
  // ??????????? 
   reg res; 
 
// module RStrigger � ???????? ? RS-???????? ?? ?-??,  
// ? RS-???????? ?? ???-??. 
// ??????????????, ??? ?? ?????? ?????? ?? ??? RS-???????? 
// ????????? ?????????? ????????. 
// ????????? ???????? ????????, ???? 
// ????????? ???????? ?????????? x ??? xdop.  
   always @(xdop or x) 
      begin 
 
// ???? ???????? ?? ??????????????? ?????? ?? ????? R,  
// ?? ? ??????? ????? 0:  
        if (~xdop) 
           res = 0; 
        else 
// ? ???? ???????? ?? ??????????????? ?????? ?? ????? S,  
// ?? ? ??????? ????? 1: 
          if (~x) 
           res = 1; 
      end 
// ??????????? ? ?????? ???????? ???????? ?? ?????:   
   assign out = !res; 
endmodule 
// ????? ?????? 
 
// ?????????? ???????? ?????? ??????????? ??????? ? ??? ??????????: 
       module Filter (OutResult, X, A, B, AInv, BInv); 
 
// ??????????? ??????????:    
  // ??????? ? ???????? 
 
   input   X, A, B;          //??????????? ??????, ?????????????? ??????? A ? B 
   output  OutResult, AInv, BInv;     //???????? ???? � ????????? �  
                          //??????????????? ?????? 
 
// ???????? ??????????? ??????, ??????????? ?????????? ???????? 
// ?????????????? ? ??????? NOT1 ? NOT2 
// ??????????? ?????????? ? ? ? ? ??????????? ????????  
// ?????????? AInv ? BInv ?????????????? 
   not NOT1 (AInv, A); 
   not NOT2 (BInv, B); 
 
// ???????? 4 ???? ?????? RSTrigger, ?.?. ? ??? ? ????? 4 ????????,  
// ?????????? ??????????????? ????????? ??????? ???????? ??????? ?????? 
   RStrigger call1 (out1, X, A); 
   RStrigger call2 (out2, X, B); 
   RStrigger call3 (out3, X, AInv); 
   RStrigger call4 (out4, X, BInv); 
 
//????? ??????, ???????????? ?????????? ???????? ? ? ?????? AND1: 
   and  AND1 (OutResult, out1, out2, out3, out4); 
endmodule 