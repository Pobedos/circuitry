LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY lab10_8 IS
	PORT
	(JK :IN STD_LOGIC;
	C :IN STD_LOGIC;
	R :IN STD_LOGIC;
	Q0 :INOUT STD_LOGIC;
	Q1 :INOUT STD_LOGIC;
	Q2 :INOUT STD_LOGIC;
	Q3 :INOUT STD_LOGIC);
END lab10_8;

ARCHITECTURE behav OF lab10_8 IS
SIGNAL P0, P1, P2, P3: STD_LOGIC;
BEGIN
Q0<=P0;
Q1<=P1;
Q2<=P2;
Q3<=P3;
process(JK, C, R, Q1, Q2, Q3, Q0)begin
	if(R='0') then
		P0<='0';
	elsif(C'event and C='1') then
		if(JK='1') then
			P0<=not(P0);
		end if;
	end if;

	if(R='0') then
		P1<='0';
	elsif(Q0'event and Q0='0') then
		if(JK='1') then
			P1<=not(P1);
		end if;
	end if;
	
	if(R='0') then
		P2<='0';
	elsif(Q1'event and Q1='0') then
		if(JK='1') then
			P2<=not(P2);
		end if;
	end if;
	
	if(R='0') then
		P3<='0';
	elsif(Q2'event and Q2='0') then
		if(JK='1') then
			P3<=not(P3);
		end if;
	end if;
	end process;
END behav;
