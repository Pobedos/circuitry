library verilog;
use verilog.vl_types.all;
entity timer_tb is
end timer_tb;
