LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fbuffer IS

	PORT
	(
		DATA0 : IN STD_LOGIC;
		DATA1 : IN STD_LOGIC;
		DATA2 : IN STD_LOGIC;
		DATA3 : IN STD_LOGIC;
		DATA4 : IN STD_LOGIC;
		DATA5 : IN STD_LOGIC;
		DATA6 : IN STD_LOGIC;
		DATA7 : IN STD_LOGIC;

		RD : IN STD_LOGIC;
		WR : IN STD_LOGIC;

		ARD0 : IN STD_LOGIC;
		ARD1 : IN STD_LOGIC;
		ARD2 : IN STD_LOGIC;

		AWR0 : IN STD_LOGIC;
		AWR1 : IN STD_LOGIC;
		AWR2 : IN STD_LOGIC;

		Q0 : INOUT STD_LOGIC;
		Q1 : INOUT STD_LOGIC;
		Q2 : INOUT STD_LOGIC;
		Q3 : INOUT STD_LOGIC;
		Q4 : INOUT STD_LOGIC;
		Q5 : INOUT STD_LOGIC;
		Q6 : INOUT STD_LOGIC;
		Q7 : INOUT STD_LOGIC;


		TMP_F0 : INOUT STD_LOGIC;
		TMP_F1 : INOUT STD_LOGIC;
		TMP_F2 : INOUT STD_LOGIC;
		TMP_F3 : INOUT STD_LOGIC;
		TMP_F4 : INOUT STD_LOGIC;
		TMP_F5 : INOUT STD_LOGIC;
		TMP_F6 : INOUT STD_LOGIC;
		TMP_F7 : INOUT STD_LOGIC;

		TMP_DFFQ00 : INOUT STD_LOGIC;
		TMP_DFFQ01 : INOUT STD_LOGIC;
		TMP_DFFQ02 : INOUT STD_LOGIC;
		TMP_DFFQ03 : INOUT STD_LOGIC;
		TMP_DFFQ04 : INOUT STD_LOGIC;
		TMP_DFFQ05 : INOUT STD_LOGIC;
		TMP_DFFQ06 : INOUT STD_LOGIC;
		TMP_DFFQ07 : INOUT STD_LOGIC;
	
		TMP_DFFQ10 : INOUT STD_LOGIC;
		TMP_DFFQ11 : INOUT STD_LOGIC;
		TMP_DFFQ12 : INOUT STD_LOGIC;
		TMP_DFFQ13 : INOUT STD_LOGIC;
		TMP_DFFQ14 : INOUT STD_LOGIC;
		TMP_DFFQ15 : INOUT STD_LOGIC;
		TMP_DFFQ16 : INOUT STD_LOGIC;
		TMP_DFFQ17 : INOUT STD_LOGIC;

		TMP_DFFQ20 : INOUT STD_LOGIC;
		TMP_DFFQ21 : INOUT STD_LOGIC;
		TMP_DFFQ22 : INOUT STD_LOGIC;
		TMP_DFFQ23 : INOUT STD_LOGIC;
		TMP_DFFQ24 : INOUT STD_LOGIC;
		TMP_DFFQ25 : INOUT STD_LOGIC;
		TMP_DFFQ26 : INOUT STD_LOGIC;
		TMP_DFFQ27 : INOUT STD_LOGIC;
	
		TMP_DFFQ30 : INOUT STD_LOGIC;
		TMP_DFFQ31 : INOUT STD_LOGIC;
		TMP_DFFQ32 : INOUT STD_LOGIC;
		TMP_DFFQ33 : INOUT STD_LOGIC;
		TMP_DFFQ34 : INOUT STD_LOGIC;
		TMP_DFFQ35 : INOUT STD_LOGIC;
		TMP_DFFQ36 : INOUT STD_LOGIC;
		TMP_DFFQ37 : INOUT STD_LOGIC;

		TMP_DFFQ40 : INOUT STD_LOGIC;
		TMP_DFFQ41 : INOUT STD_LOGIC;
		TMP_DFFQ42 : INOUT STD_LOGIC;
		TMP_DFFQ43 : INOUT STD_LOGIC;
		TMP_DFFQ44 : INOUT STD_LOGIC;
		TMP_DFFQ45 : INOUT STD_LOGIC;
		TMP_DFFQ46 : INOUT STD_LOGIC;
		TMP_DFFQ47 : INOUT STD_LOGIC;
	
		TMP_DFFQ50 : INOUT STD_LOGIC;
		TMP_DFFQ51 : INOUT STD_LOGIC;
		TMP_DFFQ52 : INOUT STD_LOGIC;
		TMP_DFFQ53 : INOUT STD_LOGIC;
		TMP_DFFQ54 : INOUT STD_LOGIC;
		TMP_DFFQ55 : INOUT STD_LOGIC;
		TMP_DFFQ56 : INOUT STD_LOGIC;
		TMP_DFFQ57 : INOUT STD_LOGIC;

		TMP_DFFQ60 : INOUT STD_LOGIC;
		TMP_DFFQ61 : INOUT STD_LOGIC;
		TMP_DFFQ62 : INOUT STD_LOGIC;
		TMP_DFFQ63 : INOUT STD_LOGIC;
		TMP_DFFQ64 : INOUT STD_LOGIC;
		TMP_DFFQ65 : INOUT STD_LOGIC;
		TMP_DFFQ66 : INOUT STD_LOGIC;
		TMP_DFFQ67 : INOUT STD_LOGIC;
	
		TMP_DFFQ70 : INOUT STD_LOGIC;
		TMP_DFFQ71 : INOUT STD_LOGIC;
		TMP_DFFQ72 : INOUT STD_LOGIC;
		TMP_DFFQ73 : INOUT STD_LOGIC;
		TMP_DFFQ74 : INOUT STD_LOGIC;
		TMP_DFFQ75 : INOUT STD_LOGIC;
		TMP_DFFQ76 : INOUT STD_LOGIC;
		TMP_DFFQ77 : INOUT STD_LOGIC;

		TMP_MUXQ0  : INOUT STD_LOGIC;
		TMP_MUXQ1  : INOUT STD_LOGIC;
		TMP_MUXQ2  : INOUT STD_LOGIC;
		TMP_MUXQ3  : INOUT STD_LOGIC;
		TMP_MUXQ4  : INOUT STD_LOGIC;
		TMP_MUXQ5  : INOUT STD_LOGIC;
		TMP_MUXQ6  : INOUT STD_LOGIC;
		TMP_MUXQ7  : INOUT STD_LOGIC
	);
	
END fbuffer;

ARCHITECTURE arch OF fbuffer IS

COMPONENT mem8
PORT( 
	  CLK	:	IN	STD_LOGIC;
	  D0	:	IN	STD_LOGIC;
      D1	:	IN	STD_LOGIC;
      D2	:	IN	STD_LOGIC;
      D3	:	IN	STD_LOGIC;
      D4	:	IN	STD_LOGIC;
      D5	:	IN	STD_LOGIC;
      D6	:	IN	STD_LOGIC;
      D7	:	IN	STD_LOGIC;

	  Q0	:	INOUT	STD_LOGIC;
      Q1	:	INOUT	STD_LOGIC;
      Q2	:	INOUT	STD_LOGIC;
      Q3	:	INOUT	STD_LOGIC;
      Q4	:	INOUT	STD_LOGIC;
      Q5	:	INOUT	STD_LOGIC;
      Q6	:	INOUT	STD_LOGIC;
      Q7	:	INOUT	STD_LOGIC
);
END COMPONENT;

COMPONENT demux8
PORT(
	E : IN STD_LOGIC;
	ADR0 : IN STD_LOGIC;
	ADR1 : IN STD_LOGIC;
	ADR2 : IN STD_LOGIC;

	F0 : INOUT STD_LOGIC;
	F1 : INOUT STD_LOGIC;
	F2 : INOUT STD_LOGIC;
	F3 : INOUT STD_LOGIC;
	F4 : INOUT STD_LOGIC;
	F5 : INOUT STD_LOGIC;
	F6 : INOUT STD_LOGIC;
	F7 : INOUT STD_LOGIC
);
END COMPONENT;

COMPONENT mux8x8
PORT
(
	ADR0 : IN STD_LOGIC;
	ADR1 : IN STD_LOGIC;
	ADR2 : IN STD_LOGIC;


	D00 : IN STD_LOGIC;
	D01 : IN STD_LOGIC;
	D02 : IN STD_LOGIC;
	D03 : IN STD_LOGIC;
	D04 : IN STD_LOGIC;
	D05 : IN STD_LOGIC;
	D06 : IN STD_LOGIC;
	D07 : IN STD_LOGIC;

	D10 : IN STD_LOGIC;
	D11 : IN STD_LOGIC;
	D12 : IN STD_LOGIC;
	D13 : IN STD_LOGIC;
	D14 : IN STD_LOGIC;
	D15 : IN STD_LOGIC;
	D16 : IN STD_LOGIC;
	D17 : IN STD_LOGIC;

	D20 : IN STD_LOGIC;
	D21 : IN STD_LOGIC;
	D22 : IN STD_LOGIC;
	D23 : IN STD_LOGIC;
	D24 : IN STD_LOGIC;
	D25 : IN STD_LOGIC;
	D26 : IN STD_LOGIC;
	D27 : IN STD_LOGIC;

	D30 : IN STD_LOGIC;
	D31 : IN STD_LOGIC;
	D32 : IN STD_LOGIC;
	D33 : IN STD_LOGIC;
	D34 : IN STD_LOGIC;
	D35 : IN STD_LOGIC;
	D36 : IN STD_LOGIC;
	D37 : IN STD_LOGIC;

	D40 : IN STD_LOGIC;
	D41 : IN STD_LOGIC;
	D42 : IN STD_LOGIC;
	D43 : IN STD_LOGIC;
	D44 : IN STD_LOGIC;
	D45 : IN STD_LOGIC;
	D46 : IN STD_LOGIC;
	D47 : IN STD_LOGIC;

	D50 : IN STD_LOGIC;
	D51 : IN STD_LOGIC;
	D52 : IN STD_LOGIC;
	D53 : IN STD_LOGIC;
	D54 : IN STD_LOGIC;
	D55 : IN STD_LOGIC;
	D56 : IN STD_LOGIC;
	D57 : IN STD_LOGIC;

	D60 : IN STD_LOGIC;
	D61 : IN STD_LOGIC;
	D62 : IN STD_LOGIC;
	D63 : IN STD_LOGIC;
	D64 : IN STD_LOGIC;
	D65 : IN STD_LOGIC;
	D66 : IN STD_LOGIC;
	D67 : IN STD_LOGIC;

	D70 : IN STD_LOGIC;
	D71 : IN STD_LOGIC;
	D72 : IN STD_LOGIC;
	D73 : IN STD_LOGIC;
	D74 : IN STD_LOGIC;
	D75 : IN STD_LOGIC;
	D76 : IN STD_LOGIC;
	D77 : IN STD_LOGIC;


	Q0 : INOUT STD_LOGIC;
	Q1 : INOUT STD_LOGIC;
	Q2 : INOUT STD_LOGIC;
	Q3 : INOUT STD_LOGIC;
	Q4 : INOUT STD_LOGIC;
	Q5 : INOUT STD_LOGIC;
	Q6 : INOUT STD_LOGIC;
	Q7 : INOUT STD_LOGIC
);	
END COMPONENT;

BEGIN

dm8 : demux8
PORT MAP( WR, AWR0, AWR1, AWR2, TMP_F0, TMP_F1, TMP_F2, TMP_F3, TMP_F4, TMP_F5, TMP_F6, TMP_F7 );

mem8_0 : mem8
PORT MAP( TMP_F0, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ00, TMP_DFFQ01, TMP_DFFQ02, TMP_DFFQ03, TMP_DFFQ04, TMP_DFFQ05, TMP_DFFQ06, TMP_DFFQ07 );
mem8_1 : mem8
PORT MAP( TMP_F1, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ10, TMP_DFFQ11, TMP_DFFQ12, TMP_DFFQ13, TMP_DFFQ14, TMP_DFFQ15, TMP_DFFQ16, TMP_DFFQ17 );
mem8_2 : mem8
PORT MAP( TMP_F2, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ20, TMP_DFFQ21, TMP_DFFQ22, TMP_DFFQ23, TMP_DFFQ24, TMP_DFFQ25, TMP_DFFQ26, TMP_DFFQ27 );
mem8_3 : mem8
PORT MAP( TMP_F3, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ30, TMP_DFFQ31, TMP_DFFQ32, TMP_DFFQ33, TMP_DFFQ34, TMP_DFFQ35, TMP_DFFQ36, TMP_DFFQ37 );
mem8_4 : mem8
PORT MAP( TMP_F4, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ40, TMP_DFFQ41, TMP_DFFQ42, TMP_DFFQ43, TMP_DFFQ44, TMP_DFFQ45, TMP_DFFQ46, TMP_DFFQ47 );
mem8_5 : mem8
PORT MAP( TMP_F5, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ50, TMP_DFFQ51, TMP_DFFQ52, TMP_DFFQ53, TMP_DFFQ54, TMP_DFFQ55, TMP_DFFQ56, TMP_DFFQ57 );
mem8_6 : mem8
PORT MAP( TMP_F6, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ60, TMP_DFFQ61, TMP_DFFQ62, TMP_DFFQ63, TMP_DFFQ64, TMP_DFFQ65, TMP_DFFQ66, TMP_DFFQ67 );
mem8_7 : mem8
PORT MAP( TMP_F7, DATA0,      DATA1,      DATA2,      DATA3,      DATA4,      DATA5,      DATA6,      DATA7,
                  TMP_DFFQ70, TMP_DFFQ71, TMP_DFFQ72, TMP_DFFQ73, TMP_DFFQ74, TMP_DFFQ75, TMP_DFFQ76, TMP_DFFQ77 );

mx8x8 : mux8x8
PORT MAP( ARD0, ARD1, ARD2,
          TMP_DFFQ00, TMP_DFFQ01, TMP_DFFQ02, TMP_DFFQ03, TMP_DFFQ04, TMP_DFFQ05, TMP_DFFQ06, TMP_DFFQ07,
		  TMP_DFFQ10, TMP_DFFQ11, TMP_DFFQ12, TMP_DFFQ13, TMP_DFFQ14, TMP_DFFQ15, TMP_DFFQ16, TMP_DFFQ17,
		  TMP_DFFQ20, TMP_DFFQ21, TMP_DFFQ22, TMP_DFFQ23, TMP_DFFQ24, TMP_DFFQ25, TMP_DFFQ26, TMP_DFFQ27,
		  TMP_DFFQ30, TMP_DFFQ31, TMP_DFFQ32, TMP_DFFQ33, TMP_DFFQ34, TMP_DFFQ35, TMP_DFFQ36, TMP_DFFQ37,
		  TMP_DFFQ40, TMP_DFFQ41, TMP_DFFQ42, TMP_DFFQ43, TMP_DFFQ44, TMP_DFFQ45, TMP_DFFQ46, TMP_DFFQ47,
		  TMP_DFFQ50, TMP_DFFQ51, TMP_DFFQ52, TMP_DFFQ53, TMP_DFFQ54, TMP_DFFQ55, TMP_DFFQ56, TMP_DFFQ57,
		  TMP_DFFQ60, TMP_DFFQ61, TMP_DFFQ62, TMP_DFFQ63, TMP_DFFQ64, TMP_DFFQ65, TMP_DFFQ66, TMP_DFFQ67,
		  TMP_DFFQ70, TMP_DFFQ71, TMP_DFFQ72, TMP_DFFQ73, TMP_DFFQ74, TMP_DFFQ75, TMP_DFFQ76, TMP_DFFQ77,
		  TMP_MUXQ0,  TMP_MUXQ1,  TMP_MUXQ2,  TMP_MUXQ3,  TMP_MUXQ4,  TMP_MUXQ5,  TMP_MUXQ6,  TMP_MUXQ7   );

mem8_out : mem8
PORT MAP( RD, TMP_MUXQ0,  TMP_MUXQ1,  TMP_MUXQ2,  TMP_MUXQ3,  TMP_MUXQ4,  TMP_MUXQ5,  TMP_MUXQ6,  TMP_MUXQ7,
		      Q0,         Q1,         Q2,         Q3,         Q4,         Q5,         Q6,         Q7         );

END arch;

CONFIGURATION conf OF fbuffer IS
	FOR arch

		FOR dm8 : demux8
			USE ENTITY work.demux8(arch);
		END FOR;
		
		FOR mem8_0, mem8_1, mem8_2, mem8_3, mem8_4, mem8_5, mem8_6, mem8_7 : mem8
			USE ENTITY work.mem8(arch);
		END FOR;
		
		FOR mx8x8 : mux8x8
			USE ENTITY work.mux8x8(arch);
		END FOR;

		FOR mem8_out : mem8
			USE ENTITY work.mem8(arch);
		END FOR;

	END FOR;
END conf;
