LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY lifo IS

	PORT
	(
		DATA0 : IN STD_LOGIC;
		DATA1 : IN STD_LOGIC;
		DATA2 : IN STD_LOGIC;
		DATA3 : IN STD_LOGIC;
		DATA4 : IN STD_LOGIC;
		DATA5 : IN STD_LOGIC;
		DATA6 : IN STD_LOGIC;
		DATA7 : IN STD_LOGIC;

		RD    : IN STD_LOGIC;
		WR    : IN STD_LOGIC;
		RESET : IN STD_LOGIC;

		Q0 : INOUT STD_LOGIC;
		Q1 : INOUT STD_LOGIC;
		Q2 : INOUT STD_LOGIC;
		Q3 : INOUT STD_LOGIC;
		Q4 : INOUT STD_LOGIC;
		Q5 : INOUT STD_LOGIC;
		Q6 : INOUT STD_LOGIC;
		Q7 : INOUT STD_LOGIC;

		FULL  : INOUT STD_LOGIC;
		EMPTY : INOUT STD_LOGIC;


		TMP_AWR0 : INOUT STD_LOGIC;
		TMP_AWR1 : INOUT STD_LOGIC;
		TMP_AWR2 : INOUT STD_LOGIC;

		TMP_ARD0 : INOUT STD_LOGIC;
		TMP_ARD1 : INOUT STD_LOGIC;
		TMP_ARD2 : INOUT STD_LOGIC;

		TMP_REQW : INOUT STD_LOGIC;
		TMP_T : INOUT STD_LOGIC;
		TMP_TI : INOUT STD_LOGIC
);
	
END lifo;

ARCHITECTURE arch OF lifo IS

COMPONENT aa5and2
PORT
(
	A		: IN	STD_LOGIC;
	B		: IN	STD_LOGIC;
	Q		: INOUT	STD_LOGIC
);
END COMPONENT;

COMPONENT rstrigger
PORT
(
	S	: IN	STD_LOGIC;
	R   : IN	STD_LOGIC;
	Q	: INOUT	STD_LOGIC;
	QI	: INOUT	STD_LOGIC
);
END COMPONENT;

COMPONENT counter
PORT
(
	CLK		:  IN	  STD_LOGIC;
	RESET	:  IN	  STD_LOGIC;
	Q1		:  INOUT  STD_LOGIC;
	Q2		:  INOUT  STD_LOGIC;
	Q3		:  INOUT  STD_LOGIC
);
END COMPONENT;

COMPONENT comp3
PORT
(
	A0 : IN STD_LOGIC;
	A1 : IN STD_LOGIC;
	A2 : IN STD_LOGIC;

	B0 : IN STD_LOGIC;
	B1 : IN STD_LOGIC;
	B2 : IN STD_LOGIC;

	AEQB : INOUT STD_LOGIC
);
END COMPONENT;

COMPONENT lbuffer
PORT
(
	DATA0 : IN STD_LOGIC;
	DATA1 : IN STD_LOGIC;
	DATA2 : IN STD_LOGIC;
	DATA3 : IN STD_LOGIC;
	DATA4 : IN STD_LOGIC;
	DATA5 : IN STD_LOGIC;
	DATA6 : IN STD_LOGIC;
	DATA7 : IN STD_LOGIC;

	RD : IN STD_LOGIC;
	WR : IN STD_LOGIC;

	Q0 : INOUT STD_LOGIC;
	Q1 : INOUT STD_LOGIC;
	Q2 : INOUT STD_LOGIC;
	Q3 : INOUT STD_LOGIC;
	Q4 : INOUT STD_LOGIC;
	Q5 : INOUT STD_LOGIC;
	Q6 : INOUT STD_LOGIC;
	Q7 : INOUT STD_LOGIC
);
END COMPONENT;


BEGIN

rcntr : counter
PORT MAP( RD, RESET, TMP_ARD0, TMP_ARD1, TMP_ARD2 );
wcntr : counter
PORT MAP( WR, RESET, TMP_AWR0, TMP_AWR1, TMP_AWR2 );
rstr : rstrigger
PORT MAP( WR, RD, TMP_T, TMP_TI );
cmp : comp3
PORT MAP( TMP_ARD0, TMP_ARD1, TMP_ARD2, TMP_AWR0, TMP_AWR1, TMP_AWR2, TMP_REQW );
fand : aa5and2
PORT MAP( TMP_T, TMP_REQW, FULL );
eand : aa5and2
PORT MAP( TMP_TI, TMP_REQW, EMPTY );
buf : lbuffer
PORT MAP( DATA0, DATA1, DATA2, DATA3, DATA4, DATA5, DATA6, DATA7, 
          RD, WR, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7 );

END arch;

CONFIGURATION conf OF lifo IS
	FOR arch

		FOR rstr : rstrigger
			USE ENTITY work.rstrigger(arch);
		END FOR;
		
		FOR rcntr, wcntr : counter
			USE ENTITY work.counter(arch);
		END FOR;

		FOR cmp : comp3
			USE ENTITY work.comp3(arch);
		END FOR;

		FOR fand, eand : aa5and2
			USE ENTITY work.aa5and2(arch);
		END FOR;

		FOR buf : lbuffer
			USE ENTITY work.lbuffer(arch);
		END FOR;

	END FOR;
END conf;

