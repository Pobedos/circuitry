LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux8x8 IS

	PORT
	(
		ADR0 : IN STD_LOGIC;
		ADR1 : IN STD_LOGIC;
		ADR2 : IN STD_LOGIC;


		D00 : IN STD_LOGIC;
		D01 : IN STD_LOGIC;
		D02 : IN STD_LOGIC;
		D03 : IN STD_LOGIC;
		D04 : IN STD_LOGIC;
		D05 : IN STD_LOGIC;
		D06 : IN STD_LOGIC;
		D07 : IN STD_LOGIC;

		D10 : IN STD_LOGIC;
		D11 : IN STD_LOGIC;
		D12 : IN STD_LOGIC;
		D13 : IN STD_LOGIC;
		D14 : IN STD_LOGIC;
		D15 : IN STD_LOGIC;
		D16 : IN STD_LOGIC;
		D17 : IN STD_LOGIC;

		D20 : IN STD_LOGIC;
		D21 : IN STD_LOGIC;
		D22 : IN STD_LOGIC;
		D23 : IN STD_LOGIC;
		D24 : IN STD_LOGIC;
		D25 : IN STD_LOGIC;
		D26 : IN STD_LOGIC;
		D27 : IN STD_LOGIC;

		D30 : IN STD_LOGIC;
		D31 : IN STD_LOGIC;
		D32 : IN STD_LOGIC;
		D33 : IN STD_LOGIC;
		D34 : IN STD_LOGIC;
		D35 : IN STD_LOGIC;
		D36 : IN STD_LOGIC;
		D37 : IN STD_LOGIC;

		D40 : IN STD_LOGIC;
		D41 : IN STD_LOGIC;
		D42 : IN STD_LOGIC;
		D43 : IN STD_LOGIC;
		D44 : IN STD_LOGIC;
		D45 : IN STD_LOGIC;
		D46 : IN STD_LOGIC;
		D47 : IN STD_LOGIC;

		D50 : IN STD_LOGIC;
		D51 : IN STD_LOGIC;
		D52 : IN STD_LOGIC;
		D53 : IN STD_LOGIC;
		D54 : IN STD_LOGIC;
		D55 : IN STD_LOGIC;
		D56 : IN STD_LOGIC;
		D57 : IN STD_LOGIC;

		D60 : IN STD_LOGIC;
		D61 : IN STD_LOGIC;
		D62 : IN STD_LOGIC;
		D63 : IN STD_LOGIC;
		D64 : IN STD_LOGIC;
		D65 : IN STD_LOGIC;
		D66 : IN STD_LOGIC;
		D67 : IN STD_LOGIC;

		D70 : IN STD_LOGIC;
		D71 : IN STD_LOGIC;
		D72 : IN STD_LOGIC;
		D73 : IN STD_LOGIC;
		D74 : IN STD_LOGIC;
		D75 : IN STD_LOGIC;
		D76 : IN STD_LOGIC;
		D77 : IN STD_LOGIC;


		Q0 : INOUT STD_LOGIC;
		Q1 : INOUT STD_LOGIC;
		Q2 : INOUT STD_LOGIC;
		Q3 : INOUT STD_LOGIC;
		Q4 : INOUT STD_LOGIC;
		Q5 : INOUT STD_LOGIC;
		Q6 : INOUT STD_LOGIC;
		Q7 : INOUT STD_LOGIC
	);
	
END mux8x8;

ARCHITECTURE arch OF mux8x8 IS

	SIGNAL Q0S, Q1S, Q2S, Q3S, Q4S, Q5S, Q6S, Q7S	: STD_LOGIC;
	
BEGIN

	PROCESS ( ADR0, ADR1, ADR2, 
              D00, D01, D02, D03, D04, D05, D06, D07,
			  D10, D11, D12, D13, D14, D15, D16, D17,
			  D20, D21, D22, D23, D24, D25, D26, D27,
			  D30, D31, D32, D33, D34, D35, D36, D37,
              D40, D41, D42, D43, D44, D45, D46, D47,
			  D50, D51, D52, D53, D54, D55, D56, D57,
			  D60, D61, D62, D63, D64, D65, D66, D67,
			  D70, D71, D72, D73, D74, D75, D76, D77 )
	BEGIN
		IF ( ADR0 = '0' AND ADR1 = '0' AND ADR2 = '0' ) THEN
			Q0S <= D00; Q1S <= D01; Q2S <= D02; Q3S <= D03; Q4S <= D04; Q5S <= D05; Q6S <= D06; Q7S <= D07;
		ELSIF ( ADR0 = '1' AND ADR1 = '0' AND ADR2 = '0' ) THEN
			Q0S <= D10; Q1S <= D11; Q2S <= D12; Q3S <= D13; Q4S <= D14; Q5S <= D15; Q6S <= D16; Q7S <= D17;
		ELSIF ( ADR0 = '0' AND ADR1 = '1' AND ADR2 = '0' ) THEN
			Q0S <= D20; Q1S <= D21; Q2S <= D22; Q3S <= D23; Q4S <= D24; Q5S <= D25; Q6S <= D26; Q7S <= D27;
		ELSIF ( ADR0 = '1' AND ADR1 = '1' AND ADR2 = '0' ) THEN
			Q0S <= D30; Q1S <= D31; Q2S <= D32; Q3S <= D33; Q4S <= D34; Q5S <= D35; Q6S <= D36; Q7S <= D37;
		ELSIF ( ADR0 = '0' AND ADR1 = '0' AND ADR2 = '1' ) THEN
			Q0S <= D40; Q1S <= D41; Q2S <= D42; Q3S <= D43; Q4S <= D44; Q5S <= D45; Q6S <= D46; Q7S <= D47;
		ELSIF ( ADR0 = '1' AND ADR1 = '0' AND ADR2 = '1' ) THEN
			Q0S <= D50; Q1S <= D51; Q2S <= D52; Q3S <= D53; Q4S <= D54; Q5S <= D55; Q6S <= D56; Q7S <= D57;
		ELSIF ( ADR0 = '0' AND ADR1 = '1' AND ADR2 = '1' ) THEN
			Q0S <= D60; Q1S <= D61; Q2S <= D62; Q3S <= D63; Q4S <= D64; Q5S <= D65; Q6S <= D66; Q7S <= D67;
		ELSIF ( ADR0 = '1' AND ADR1 = '1' AND ADR2 = '1' ) THEN
			Q0S <= D70; Q1S <= D71; Q2S <= D72; Q3S <= D73; Q4S <= D74; Q5S <= D75; Q6S <= D76; Q7S <= D77;
		END IF;
	END PROCESS;

	Q0 <= Q0S; Q1 <= Q1S; Q2 <= Q2S; Q3 <= Q3S;
	Q4 <= Q4S; Q5 <= Q5S; Q6 <= Q6S; Q7 <= Q7S;

END arch;
