LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mem8x8 IS
PORT( CLK	:	IN	STD_LOGIC;
	  D0	:	IN	STD_LOGIC;
      D1	:	IN	STD_LOGIC;
      D2	:	IN	STD_LOGIC;
      D3	:	IN	STD_LOGIC;
      D4	:	IN	STD_LOGIC;
      D5	:	IN	STD_LOGIC;
      D6	:	IN	STD_LOGIC;
      D7	:	IN	STD_LOGIC;

	  T0Q0	:	INOUT	STD_LOGIC;
      T0Q1	:	INOUT	STD_LOGIC;
      T0Q2	:	INOUT	STD_LOGIC;
      T0Q3	:	INOUT	STD_LOGIC;
      T0Q4	:	INOUT	STD_LOGIC;
      T0Q5	:	INOUT	STD_LOGIC;
      T0Q6	:	INOUT	STD_LOGIC;
      T0Q7	:	INOUT	STD_LOGIC;	

	  T1Q0	:	INOUT	STD_LOGIC;
      T1Q1	:	INOUT	STD_LOGIC;
      T1Q2	:	INOUT	STD_LOGIC;
      T1Q3	:	INOUT	STD_LOGIC;
      T1Q4	:	INOUT	STD_LOGIC;
      T1Q5	:	INOUT	STD_LOGIC;
      T1Q6	:	INOUT	STD_LOGIC;
      T1Q7	:	INOUT	STD_LOGIC;	

	  T2Q0	:	INOUT	STD_LOGIC;
      T2Q1	:	INOUT	STD_LOGIC;
      T2Q2	:	INOUT	STD_LOGIC;
      T2Q3	:	INOUT	STD_LOGIC;
      T2Q4	:	INOUT	STD_LOGIC;
      T2Q5	:	INOUT	STD_LOGIC;
      T2Q6	:	INOUT	STD_LOGIC;
      T2Q7	:	INOUT	STD_LOGIC;	

	  T3Q0	:	INOUT	STD_LOGIC;
      T3Q1	:	INOUT	STD_LOGIC;
      T3Q2	:	INOUT	STD_LOGIC;
      T3Q3	:	INOUT	STD_LOGIC;
      T3Q4	:	INOUT	STD_LOGIC;
      T3Q5	:	INOUT	STD_LOGIC;
      T3Q6	:	INOUT	STD_LOGIC;
      T3Q7	:	INOUT	STD_LOGIC;	

	  T4Q0	:	INOUT	STD_LOGIC;
      T4Q1	:	INOUT	STD_LOGIC;
      T4Q2	:	INOUT	STD_LOGIC;
      T4Q3	:	INOUT	STD_LOGIC;
      T4Q4	:	INOUT	STD_LOGIC;
      T4Q5	:	INOUT	STD_LOGIC;
      T4Q6	:	INOUT	STD_LOGIC;
      T4Q7	:	INOUT	STD_LOGIC;	

	  T5Q0	:	INOUT	STD_LOGIC;
      T5Q1	:	INOUT	STD_LOGIC;
      T5Q2	:	INOUT	STD_LOGIC;
      T5Q3	:	INOUT	STD_LOGIC;
      T5Q4	:	INOUT	STD_LOGIC;
      T5Q5	:	INOUT	STD_LOGIC;
      T5Q6	:	INOUT	STD_LOGIC;
      T5Q7	:	INOUT	STD_LOGIC;	

	  T6Q0	:	INOUT	STD_LOGIC;
      T6Q1	:	INOUT	STD_LOGIC;
      T6Q2	:	INOUT	STD_LOGIC;
      T6Q3	:	INOUT	STD_LOGIC;
      T6Q4	:	INOUT	STD_LOGIC;
      T6Q5	:	INOUT	STD_LOGIC;
      T6Q6	:	INOUT	STD_LOGIC;
      T6Q7	:	INOUT	STD_LOGIC;	

	  Q0	:	INOUT	STD_LOGIC;
      Q1	:	INOUT	STD_LOGIC;
      Q2	:	INOUT	STD_LOGIC;
      Q3	:	INOUT	STD_LOGIC;
      Q4	:	INOUT	STD_LOGIC;
      Q5	:	INOUT	STD_LOGIC;
      Q6	:	INOUT	STD_LOGIC;
      Q7	:	INOUT	STD_LOGIC
);
END mem8x8;

ARCHITECTURE arch OF mem8x8 IS

COMPONENT mem8
PORT( 
	  CLK	:	IN	STD_LOGIC;
	  D0	:	IN	STD_LOGIC;
      D1	:	IN	STD_LOGIC;
      D2	:	IN	STD_LOGIC;
      D3	:	IN	STD_LOGIC;
      D4	:	IN	STD_LOGIC;
      D5	:	IN	STD_LOGIC;
      D6	:	IN	STD_LOGIC;
      D7	:	IN	STD_LOGIC;

	  Q0	:	INOUT	STD_LOGIC;
      Q1	:	INOUT	STD_LOGIC;
      Q2	:	INOUT	STD_LOGIC;
      Q3	:	INOUT	STD_LOGIC;
      Q4	:	INOUT	STD_LOGIC;
      Q5	:	INOUT	STD_LOGIC;
      Q6	:	INOUT	STD_LOGIC;
      Q7	:	INOUT	STD_LOGIC
);
END COMPONENT;

BEGIN

mm0 : mem8
PORT MAP ( CLK, D0, D1, D2, D3, D4, D5, D6, D7, T0Q0, T0Q1, T0Q2, T0Q3, T0Q4, T0Q5, T0Q6, T0Q7 );
mm1 : mem8
PORT MAP ( CLK, T0Q0, T0Q1, T0Q2, T0Q3, T0Q4, T0Q5, T0Q6, T0Q7, T1Q0, T1Q1, T1Q2, T1Q3, T1Q4, T1Q5, T1Q6, T1Q7 );
mm2 : mem8
PORT MAP ( CLK, T1Q0, T1Q1, T1Q2, T1Q3, T1Q4, T1Q5, T1Q6, T1Q7, T2Q0, T2Q1, T2Q2, T2Q3, T2Q4, T2Q5, T2Q6, T2Q7 );
mm3 : mem8
PORT MAP ( CLK, T2Q0, T2Q1, T2Q2, T2Q3, T2Q4, T2Q5, T2Q6, T2Q7, T3Q0, T3Q1, T3Q2, T3Q3, T3Q4, T3Q5, T3Q6, T3Q7 );
mm4 : mem8
PORT MAP ( CLK, T3Q0, T3Q1, T3Q2, T3Q3, T3Q4, T3Q5, T3Q6, T3Q7, T4Q0, T4Q1, T4Q2, T4Q3, T4Q4, T4Q5, T4Q6, T4Q7 );
mm5 : mem8
PORT MAP ( CLK, T4Q0, T4Q1, T4Q2, T4Q3, T4Q4, T4Q5, T4Q6, T4Q7, T5Q0, T5Q1, T5Q2, T5Q3, T5Q4, T5Q5, T5Q6, T5Q7 );
mm6 : mem8
PORT MAP ( CLK, T5Q0, T5Q1, T5Q2, T5Q3, T5Q4, T5Q5, T5Q6, T5Q7, T6Q0, T6Q1, T6Q2, T6Q3, T6Q4, T6Q5, T6Q6, T6Q7 );
mm7 : mem8
PORT MAP ( CLK, T6Q0, T6Q1, T6Q2, T6Q3, T6Q4, T6Q5, T6Q6, T6Q7, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7 );

END arch;

CONFIGURATION conf OF mem8x8 IS
	FOR arch

		FOR mm0, mm1, mm2, mm3, mm4, mm5, mm6, mm7 : mem8
			USE ENTITY work.mem8 (arch);
		END FOR;

	END FOR;
END conf;

