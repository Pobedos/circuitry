library ieee;
use ieee.std_logic_1164.all;

package row_type is
    type row is array (0 to 3) of integer;
end package;

